module ripple_carry_adder (in0, in1, out, cout,s_overflow,u_overflow);
// declare input signals
input [3:0] in0;
input [3:0] in1;

// declare output signals
output [3:0] out;
output cout;
output s_overflow;
output u_overflow;

// here is your design

endmodule




