// ===================================================// 
//  Question 2  4-bit Ping_Pong_Counter     	      //
// ===================================================//

module Ping_Pong_Counter (CLK, RESET_n, enable, direction, out);
	
	input CLK, RESET_n;
	input enable;
	output direction;
	output [4-1:0] out;

endmodule
